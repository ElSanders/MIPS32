library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity DataMemory is
	Port( CLK, WRITE_ENABLE, READ_ENABLE: in STD_LOGIC := '0';
			ENABLE: in STD_LOGIC :='0';
			RW_ADDRESS,WRITE_DATA: in STD_LOGIC_VECTOR(31 downto 0):="00000000000000000000000000000000";
		   READ_DATA: out STD_LOGIC_VECTOR(31 downto 0):="00000000000000000000000000000000"
		  );
end DataMemory;

architecture Behavioral of DataMemory is

begin

PROCESS (RW_ADDRESS,ENABLE,WRITE_ENABLE,READ_ENABLE,CLK)
	SUBTYPE REGISTRO IS STD_LOGIC_VECTOR (31 DOWNTO 0);
		TYPE REG_BANK IS ARRAY (0 TO 31) OF REGISTRO;
		VARIABLE DATA_MEMORY: REG_BANK := (
													"00000000000000000000000000000001",
													"00000000000000000000000000000010",
													"00000000000000000000000000000011",
													"00000000000000000000000000000100",
													"00000000000000000000000000000101",
													"00000000000000000000000000000111",
													"00000000000000000000000000001000",
													"00000000000000000000000000001001",
													OTHERS => (OTHERS => '0')
		 );
		 VARIABLE ADDRESS: INTEGER;
	BEGIN
	 IF( ENABLE = '1')THEN
	 IF (READ_ENABLE = '1' and WRITE_ENABLE = '0') THEN
		ADDRESS:= TO_INTEGER(UNSIGNED(RW_ADDRESS(6 downto 2)));
		READ_DATA <= DATA_MEMORY(ADDRESS);
		ELSIF (WRITE_ENABLE = '1' and READ_ENABLE = '0' and CLK='0' and CLK'EVENT) THEN
			 ADDRESS:= TO_INTEGER(UNSIGNED(RW_ADDRESS(6 downto 2)));
			 READ_DATA <= "00000000000000000000000000000000";
			 DATA_MEMORY(ADDRESS):= WRITE_DATA;
	 ELSE NULL;
	 END IF;
ELSE NULL;
END IF;
END PROCESS;


end Behavioral;

